module hwtb();
   
endmodule : hwtb