module HDMI_Controller
  (
   input bit 	     clk,
   output bit 	     vsync, hsync,
   output bit [31:0] color
   );
   
   
endmodule : HDMI_Controller