 
module ASCII2Bitmap
   (input logic  [7:0]  char,
    output logic [149:0]     bitmap);

    always_comb begin
      case (char)
	// 0 := 48 [0x30]
	8'h30 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6DB7FFFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB6DB7FFFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 1 := 49 [0x31]
	8'h31 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFEDB7FFFFFEC937FFFFFEC937FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 2 := 50 [0x32]
	8'h32 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFEDB7EDB7FFFFFFEDB7FFFFFEDB7FFFFEC937FFFFEC937FFFFFEDB7FFFFFEC8000137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 3 := 51 [0x33]
	8'h33 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC80137FFFEDB6C937FFFFFEC937FFFFEC937FFFFFFEC937FFFFFFEDB7FFEDB7EDB7FFEDB6C937FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 4 := 52 [0x34]
	8'h34 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFEDB7FFFFFEC937FFFFFEC937FFFFEDA5B7FFFEDB6DB7FFFEDB6DB7FFEC8000137FFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 5 := 53 [0x35]
	8'h35 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC800137FFEDB7FFFFFFEDB7FFFFFFEC80137FFFEDB6C937FFFFFFEDB7FFFFFFEDB7FFEDB6C937FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 6 := 54 [0x36]
	8'h36 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFEDB7FFFFFFEC80137FFFEDB6C937FFEDB7EDB7FFEDB7EDB7FFEDB6C937FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 7 := 55 [0x37]
	8'h37 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC800137FFFFFFEDB7FFFFFEDB7FFFFFFEDB7FFFFFEDB7FFFFFFEDB7FFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 8 := 56 [0x38]
	8'h38 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFEDB6C937FFFEC8137FFFEDB6C937FFEDB7EDB7FFEDB7EDB7FFEDB6C937FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// 9 := 57 [0x39]
	8'h39 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFEDB7EDB7FFEDB7EDB7FFEDB6C937FFFEC925B7FFFFFFEDB7FFEDB6DB7FFFFEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// A := 65 [0x41]
	8'h41 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFEC937FFFFFEC937FFFFEC80137FFFEDB6DB7FFFEDB6DB7FFEC8000137FEDB7FEDB7FEDB7FEDB7EC937FEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// B := 66 [0x42]
	8'h42 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC800137FFEDB7EC937FEDB7FEDB7FEDB7FEDB7FEC800137FFEDB7FEDB7FEDB7FEDB7FEDB7FEDB7FEC800137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// C := 67 [0x43]
	8'h43 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFEC8137FFFEDB7EDB7FEDB7FFEDB7EDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFEDB7FEDB7EDB7FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// D := 68 [0x44]
	8'h44 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC800137FFEDB7FEDB7FEDB7FEC937EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FEC937EDB7FEDB7FEC800137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// E := 69 [0x45]
	8'h45 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC8000137FEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEC8000137FEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEC8000137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// F := 70 [0x46]
	8'h46 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC8000137FEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEC800137FFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// G := 71 [0x47]
	8'h47 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFEC80137FFEDB7EC937EDB7FFEDB7EDB7FFFFFFEDB7EC8137EDB7FFEC936DB7FFEC937EDB7EC8137FEC8136DB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// H := 72 [0x48]
	8'h48 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EC80000137EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// I := 73 [0x49]
	8'h49 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// J := 74 [0x4A]
	8'h4A : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFEDB7EDB7FFEC936DB7FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// K := 75 [0x4B]
	8'h4B : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FEDB7FEDB7EDB7FFEDB6DB7FFFEDA4937FFFEC80137FFFEDB6C937FFEDB7EDB7FFEDB7FEDB7FEDB7FEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// L := 76 [0x4C]
	8'h4C : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEC800137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// M := 77 [0x4D]
	8'h4D : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC937FEC936C937FEC936C937FEC936DA5B6DA5B6DA5B6DA5B6DA5B6DA5B6DB6C936DB6DB6C936DB6DB6C936DB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// N := 78 [0x4E]
	8'h4E : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFEDB7EC937FEDB7EC8137EDB7EDA5B7EDB7EDB6DB6DB7EDB6C925B7EDB7EDA5B7EDB7FEC937EDB7FEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// O := 79 [0x4F]
	8'h4F : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFEC80137FEC937EC937EDB7FFEDB7EDB7FFFEDA4937FFFEDB6DB7FFFEDB6DB7FFEDB7EC937EC937FFEC80137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// P := 80 [0x50]
	8'h50 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC800137FFEDB7FEDB7FEDB7FEDB7FEDB7FEDB7FEC8000137FEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// Q := 81 [0x51]
	8'h51 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFEC80137FEC937EC937EDB7FFEDB7EDB7FFFEDA4937FFFEDB6DB7FFFEDB6DB7FFEDB7EC937EC937FFEC800137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// R := 82 [0x52]
	8'h52 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC8000137FEDB7FEC937EDB7FFEDB7EDB7FEDB7FEC8000137FEDB7FEDB7FEDB7FEC937EDB7FFEDB7EDB7FFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// S := 83 [0x53]
	8'h53 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEC80137FFEC936C937FEDB7FEDB7FEC937FFFFFFFEC8137FFFFFFFEDB7FEDB7FEDB7FEC937EDB7FFEC80137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// T := 84 [0x54]
	8'h54 : bitmap = 150'hFFFFFFFFFFFFFFFFFEC80000137FFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// U := 85 [0x55]
	8'h55 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EC937EDB7FFEC80137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// V := 86 [0x56]
	8'h56 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FEC937EDB7FEDB7FEDB7FEDB7FFEDB6C937FFEDB6DB7FFFEDB6DB7FFFFEC8137FFFFEC937FFFFFEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// W := 87 [0x57]
	8'h57 : bitmap = 150'hFFFFFFFFFFFFFFFFFEC937EDB7FFEDB7EC937FEDB6C8137FEDB6DA5B7FEC925A4937FEDA5B6DB7FEC937EC937EC937EC937EC937FEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// X := 88 [0x58]
	8'h58 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FEDB7FEC936C937FFEDB6DB7FFFFEC937FFFFFEC937FFFFFEC937FFFFEDB6DB7FFEC936C937FEDB7FEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// Y := 89 [0x59]
	8'h59 : bitmap = 150'hFFFFFFFFFFFFFFFFFEC937FEC937EDB7FEDB7FFEDB6DB7FFFEC925B7FFFFEC937FFFFFEC937FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// Z := 90 [0x5A]
	8'h5A : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC8000137FFFFFEC937FFFFEC937FFFFFEDB7FFFFFEDB7FFFFFEC937FFFFEC937FFFFFEDB7FFFFFEC80000137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// a := 97 [0x61]
	8'h61 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFFFFEC937FFEC800137FFEDB7EDB7FFEDB6C937FFEC8125B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// b := 98 [0x62]
	8'h62 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEC80137FFFEDB6C937FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB6C937FFEC80137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// c := 99 [0x63]
	8'h63 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6DB7FFFEDB7FFFFFEDB7FFFFFFEC937FFFFFFEDB6DB7FFFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// d := 100 [0x64]
	8'h64 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFEC925B7FFEDB6C937FEC937EDB7FEDB7FEDB7FEC937EDB7FFEDB6C937FFFEC925B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// e := 101 [0x65]
	8'h65 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFEDB7EDB7FFEC800137FFEDB7FFFFFFEDB6C937FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// f := 102 [0x66]
	8'h66 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEC937FFFFFEDB7FFFFFEC8137FFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// g := 103 [0x67]
	8'h67 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC925B7FFEDB6C937FEC937EDB7FEDB7FEDB7FEC937EDB7FFEDB6C937FFFEC925B7FFFFFFEDB7FFEDB6DB7FFFFEC8137FFFFFFFFFFFF;
	// h := 104 [0x68]
	8'h68 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDA4937FFFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// i := 105 [0x69]
	8'h69 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// j := 106 [0x6A]
	8'h6A : bitmap = 150'hFFFFFFFFFFFFFFFFFFFEDB7FFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFEDB7FFFFFFFFFFFFFFF;
	// k := 107 [0x6B]
	8'h6B : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB6DB7FFFEDA5B7FFFFEC8137FFFFEC8137FFFFEDA4937FFFEDB6DB7FFFEDB6C937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// l := 108 [0x6C]
	8'h6C : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// m := 109 [0x6D]
	8'h6D : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC801248136DB6C936DB6DB6C936DB6DB6C936DB6DB6C936DB6DB6C936DB6DB6C936DB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// n := 110 [0x6E]
	8'h6E : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDA4937FFFEDB6C937FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// o := 111 [0x6F]
	8'h6F : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC8137FFFEDB6C937FFEDB7EDB7FEC937EDB7FFEDB7EDB7FFEDB6C937FFFEC8137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// p := 112 [0x70]
	8'h70 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC80137FFFEDB6C937FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB6C937FFEC80137FFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFF;
	// q := 113 [0x71]
	8'h71 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC925B7FFEDB6C937FEC937EDB7FEDB7FEDB7FEC937EDB7FFEDB6C937FFFEC925B7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFF;
	// r := 114 [0x72]
	8'h72 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDA5B7FFFFEC937FFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// s := 115 [0x73]
	8'h73 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC8137FFFFEDB6DB7FFFEDB7FFFFFFFEC937FFFFFFFEDB7FFFEDB6DB7FFFEC80137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// t := 116 [0x74]
	8'h74 : bitmap = 150'hFFFFFFFFFFFFFFFFFFEDB7FFFFFFEDB7FFFFFEC8137FFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEDB7FFFFFFEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// u := 117 [0x75]
	8'h75 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB7EDB7FFEDB6C937FFEC8125B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// v := 118 [0x76]
	8'h76 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDB7FEDB7FFEDB6DB7FFFEDB6DB7FFFEDB6DB7FFFFEC937FFFFFEC937FFFFFEC937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// w := 119 [0x77]
	8'h77 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDB7EDB6DB6C924936DB7EDA4936DB7EDA5A5A5B7EC8124937FEC936C937FFEDB6C937FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// x := 120 [0x78]
	8'h78 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDB6DB7FFFEDB6DB7FFFFEC937FFFFFEC937FFFFFEC937FFFFEDB6DB7FFFEDB6DB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
	// y := 121 [0x79]
	8'h79 : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDB7EC937FFEDB6DB7FFFEDB6DB7FFFEDB6DB7FFFFEC937FFFFFEC937FFFFFEC937FFFFFEDB7FFFFFFEDB7FFFFFEDB7FFFFFFFFFFFFFFF;
	// z := 122 [0x7A]
	8'h7A : bitmap = 150'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC80137FFFFFFEDB7FFFFFEDB7FFFFFEDB7FFFFFEC937FFFFFEDB7FFFFFEC800137FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

      endcase
    end
endmodule : ASCII2Bitmap
